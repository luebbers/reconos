--
-- \file %%%FILENAME%%%
--
-- %%%SHORT_DESCRIPTION%%%
--
-- %%%LONG_DESCRIPTION%%%
--
-- \author     %%%REALNAME%%% <%%%EMAIL%%%>
-- \date       %%%DATE%%%
--
-----------------------------------------------------------------------------
-- %%%RECONOS_COPYRIGHT_BEGIN%%%
-- %%%RECONOS_COPYRIGHT_END%%%
-----------------------------------------------------------------------------
--

