../thread.vhd