-------------------------------------------------------------------------------
-- $Id: command_fifo.vhd,v 1.1 2005/02/18 15:30:22 wirthlin Exp $
-------------------------------------------------------------------------------
-- srl_fifo.vhd
-------------------------------------------------------------------------------
--
--                  ****************************
--                  ** Copyright Xilinx, Inc. **
--                  ** All rights reserved.   **
--                  ****************************
--
-------------------------------------------------------------------------------
-- Filename:        
--
-- Description:     
--                  
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   
--              
--
-------------------------------------------------------------------------------
-- Author:          goran
-- Revision:        $Revision: 1.1 $
-- Date:            $Date: 2005/02/18 15:30:22 $
--
-- History:
--
-------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x" 
--      reset signals:                          "rst", "rst_n" 
--      generics:                               "C_*" 
--      user defined types:                     "*_TYPE" 
--      state machine next state:               "*_ns" 
--      state machine current state:            "*_cs" 
--      combinatorial signals:                  "*_com" 
--      pipelined or register delay signals:    "*_d#" 
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce" 
--      internal version of output port         "*_i"
--      device pins:                            "*_pin" 
--      ports:                                  - Names begin with Uppercase 
--      processes:                              "*_PROCESS" 
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
-------------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;

library UNISIM;
use UNISIM.all;
use UNISIM.vcomponents.all;

entity command_fifo is
  port (
    Clk         : in  std_logic;
    Reset       : in  std_logic;
    NextCommand : in  std_logic;
    CommandNum  : out std_logic_vector(8 downto 0);
    Data        : out std_logic_vector(15 downto 0);
    Address     : out std_logic_vector(6 downto 0);
    ValidCommand: out std_logic
    );
end entity command_fifo;


-- Commands for AC97:
--     WriteAC97Reg(0x0,0x0); // reset registers
--     WriteAC97Reg(0x2,0x808); // master volume (0db gain)
--     WriteAC97Reg(0xa,0x8000); // mute PC beep
--     WriteAC97Reg(0x4,0x808); // headphone vol (aux out)
--     WriteAC97Reg(0x18,0x808); // pcmoutvol (amp out line)
--     WriteAC97Reg(0x1a,0x404); // record source (line in for left and right)
--     WriteAC97Reg(0x1c,0x008); // record gain (8 steps of 1.5 dB = +12.0 dB)
--     WriteAC97Reg(0x20,0x1); // bypass 3d sound

-- 80000000
-- 80020808
-- 800a8000
-- 80040808
-- 80180808
-- 801a0404
-- 801c0008
-- 80200001

-- 80200001801c0008801a04048018080880040808800a80008002080880000000


architecture IMP of command_fifo is

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0a : string;
  attribute INIT_0b : string;
  attribute INIT_0c : string;
  attribute INIT_0d : string;
  attribute INIT_0e : string;
  attribute INIT_0f : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1a : string;
  attribute INIT_1b : string;
  attribute INIT_1c : string;
  attribute INIT_1d : string;
  attribute INIT_1e : string;
  attribute INIT_1f : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2a : string;
  attribute INIT_2b : string;
  attribute INIT_2c : string;
  attribute INIT_2d : string;
  attribute INIT_2e : string;
  attribute INIT_2f : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3a : string;
  attribute INIT_3b : string;
  attribute INIT_3c : string;
  attribute INIT_3d : string;
  attribute INIT_3e : string;
  attribute INIT_3f : string;


  attribute INIT_00 of u1 : label is
    "80200001801c0008801a04048018080880040808800a80008002080880000000";
  attribute INIT_01 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_02 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_03 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_04 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_05 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_06 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_07 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_08 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_09 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_0a of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_0b of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_0c of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_0d of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_0e of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_0f of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_10 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_11 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_12 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_13 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_14 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_15 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_16 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_17 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_18 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_19 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_1a of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_1b of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_1c of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_1d of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_1e of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_1f of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_20 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_21 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_22 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_23 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_24 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_25 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_26 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_27 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_28 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_29 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_2a of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_2b of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_2c of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_2d of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_2e of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_2f of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_30 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_31 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_32 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_33 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_34 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_35 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_36 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_37 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_38 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_39 of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_3a of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_3b of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_3c of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_3d of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_3e of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";
  attribute INIT_3f of u1 : label is
    "0000000000000000000000000000000000000000000000000000000000000000";

  component RAMB16_S36
    generic (
      INIT       : bit_vector := X"000000000";
      SRVAL      : bit_vector := X"000000000";
      write_mode : string     := "WRITE_FIRST";
  
      INITP_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_00  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F  : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      );
  
    port (
      DO   : out std_logic_vector (31 downto 0);
      DOP  : out std_logic_vector (3 downto 0);
      
      ADDR : in  std_logic_vector (8 downto 0);
      CLK  : in  std_ulogic;
      DI   : in  std_logic_vector (31 downto 0);
      DIP  : in  std_logic_vector (3 downto 0);
      EN   : in  std_ulogic;
      SSR  : in  std_ulogic;
      WE   : in  std_ulogic
      );
  
  end component;

  signal xram_di : std_logic_vector(31 downto 0);    -- BlockRAM data in (zero)
  signal command_addr : unsigned(8 downto 0);    -- BlockRAM data in (zero)
  signal xram_addr : std_logic_vector(8 downto 0);    -- BlockRAM data in (zero)
  signal xram_dip : std_logic_vector(3 downto 0);    -- BlockRAM data in (zero)
  signal xram_dop : std_logic_vector(3 downto 0);    -- BlockRAM data out
  signal xram_en : std_logic;                        -- BlockRAM enable (always on)
  signal xram_we : std_logic;                        -- BlockRAM write enable (zero)
  signal xram_reset : std_logic;                     -- BlockRAM reset (zero)
  signal xram_do : std_logic_vector(31 downto 0);
begin
  
  -- address (need to define)
  block_ram_address_PROCESS : process (Clk) is
  begin
    if Clk'event and Clk = '1' then
      if Reset = '1' then
        command_addr <= (others => '0');
      elsif NextCommand = '1' then
        command_addr <= command_addr + 1;
      end if;
    end if;
  end process;
  
  -- Define input signals to BlockRam
  xram_di <= (others => '0');           -- no data in
  xram_dip <= (others => '0');          -- 2-bit data (not used)
  xram_en <= '1';                       -- always enabled
  xram_we <= '0';                       -- do not need to write
  xram_reset <= '0';                  

  Data <= xram_do(15 downto 0);
  Address <= xram_do(22 downto 16);
  ValidCommand <= xram_do(31);
  
  -- Instance the BlockRam
  u1: RAMB16_S36
--translate_off
-- Note that the these generic map values are used for simulation
-- only. To insure that the simulation matches the actual ram values,
-- make sure that the attributes used above are the same as the
-- generics used below.
  generic map (
    INIT_00 =>
    X"80200001801c0008801a04048018080880040808800a80008002080880000000",
    INIT_01 =>
    X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0a =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0b =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0c =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0d =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0e =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0f =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_10 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1a =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1b =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1c =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1d =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1e =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1f =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2a =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2b =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2c =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2d =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2e =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2f =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3a =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3b =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3c =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3d =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3e =>
       X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3f =>
       X"0000000000000000000000000000000000000000000000000000000000000000"

  )
--translate_on
    port map(
           di => xram_di,
           dip => xram_dip,
           addr => xram_addr,
           do => xram_do,
           dop => xram_dop,
           clk => clk,
           SSR => xram_reset,
           EN => xram_en,
           WE => xram_we
         );
    xram_addr <= CONV_STD_LOGIC_VECTOR(command_addr, command_addr'length);

  CommandNum <= xram_addr;
  
end architecture IMP;
