#==========================================================================
# 
#       mouse_virtex4.cdl
# 
#       eCos configuration data for the Xilinx VIRTEX4 mouse
#       Taken from the Xilinx ML300 mouse
# 
#==========================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
#==========================================================================
######DESCRIPTIONBEGIN####
# 
# Author(s):    gthomas
# Contributors: gthomas, cduclos
# Date:         2002-03-03
#               2005-04-19                
# Purpose:      
# Description:  Mouse drivers for Xilinx VIRTEX4
# 
#####DESCRIPTIONEND####
# 
#==========================================================================

cdl_package CYGPKG_DEVS_MOUSE_VIRTEX4 {
    display     "Mouse driver for virtex4"
    include_dir cyg/io

#    active_if   CYGPKG_IO_FILEIO
#    requires    CYGPKG_IO
#    requires    CYGFUN_KERNEL_API_C
#    requires    CYGPKG_HAL_POWERPC_VIRTEX4
# CMDV: Originally this was !CYGSEM_VIRTEX4_LCD_COMM
    active_if   CYGSEM_VIRTEX4_LCD_COMM

    compile       -library=libextras.a virtex4_mouse.c

    description "Mouse driver for the Xilinx VIRTEX4"

    cdl_component CYGPKG_DEVS_MOUSE_VIRTEX4_OPTIONS {
        display "options"
        flavor  none
        no_define

        cdl_option CYGPKG_DEVS_MOUSE_VIRTEX4_CFLAGS {
            display       "Additional compiler flags"
            flavor        data
            no_define
            default_value { "" }
            description "
               This option modifies the set of compiler flags for
               building the mousescreen driver package. These flags
               are used in addition to the set of global flags."
        }

        cdl_option CYGDAT_DEVS_MOUSE_VIRTEX4_NAME {
            display "Device name for the mouse driver"
            flavor data
            default_value {"\"/dev/mouse\""}
            description " This option specifies the name of the mouse device"
        }

        cdl_option CYGNUM_DEVS_MOUSE_VIRTEX4_BUFFER_SIZE {
            display "Number of bytes the driver can buffer"
            flavor data
            default_value { 128 }
            description "
                This option defines the size of the mouse device internal
            buffer. The cyg_io_read() function will return as many of these
            as there is space for in the buffer passed."
        }
    }
}
