#====================================================================
#
#      virtex4_eth_drivers.cdl
#
#====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
## Copyright (C) 2003, 2004, 2005 Mind n.v.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Jan Olbrechts
# Original data:  
# Contributors:   
# Date:           2005-11-08
#
#####DESCRIPTIONEND####
#
#====================================================================

cdl_package MNDPKG_DEVS_ETH_POWERPC_VIRTEX4_SGDMATEMAC {
    display       "Xilinx VIRTEX4 (PPC405) gigabit ethernet support"
    description   "Efficient ethernet driver for Xilinx VIRTEX4."

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_HAL_POWERPC 
    requires      CYGPKG_HAL_POWERPC_VIRTEX4
    requires      CYGHWR_DEVS_ETH_PHY_VIRTEX4
    active_if     MNDHWR_VIRTEX4_SGDMATEMAC

    include_dir   .
    include_files ; # none _exported_ whatsoever

    implements    CYGHWR_NET_DRIVERS
    implements    CYGHWR_NET_DRIVER_ETH0

    compile       -library=libextras.a if_virtex4_temac_sgdma.c

    # Debug I/O during network stack initialization is not reliable
    requires { !CYGPKG_NET || CYGPKG_NET_FORCE_SERIAL_CONSOLE == 1 }
    cdl_component MNDPKG_DEVS_ETH_POWERPC_VIRTEX4_SGDMATEMAC_OPTIONS {
        display "MPC8xxx VIRTEX4 ethernet driver build options"
        flavor  none
	no_define

        cdl_option MNDPKG_DEVS_ETH_POWERPC_VIRTEX4_SGDMATEMAC_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS" }
            description   "
                This option modifies the set of compiler flags for
                building the MPC8xxx VIRTEX4 ethernet driver package. 
		These flags are used in addition to the set of global 
		flags."
        }
    }
}

