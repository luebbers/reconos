../../../../src/hwt_data.vhd