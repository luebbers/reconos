../../../../src/hwt_mutex.vhd